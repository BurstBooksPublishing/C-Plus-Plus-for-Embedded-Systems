module clock_gating (
input clk,
input stall_signal,
output reg gated_clk_stage2,
output reg gated_clk_stage3
);
// Your implementation here
endmodule